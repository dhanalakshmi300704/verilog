module top_module(
    output zero
);// Modulemodule top_module( 
    
endmodule
